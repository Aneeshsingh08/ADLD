module t_fsm();


