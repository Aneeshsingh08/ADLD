module t_a();
parameter n=4;

wire front,back;
wire [3:0] slot;
reg start,clk;
reg [n-1:0] pswd,vn;

park dut(front,back,slot,clk,start,pswd,vn);

always #5 clk=~clk;

initial 
 begin
  clk=1'b1;
  start=1'b0;
  pswd=4'b0000;
   vn=4'b0000;
	#10 start=1'b1;
	    vn=4'b1000;
	    pswd=4'b1001;
	 #10  pswd=4'b1010;
	 
	#10 start=1'b0;
	#10 pswd=4'b0000;
	
	#10 start=1'b1;
	    vn=4'b1100;
	
	#10 pswd=4'b1101;
	#20 pswd=4'b1010;
	#10 start=1'b0;
	
	
  end

initial 
 begin
	$monitor ($time,"Front=%2d,Back=%2d,slot=%2d",front,back,slot);
	#200  $finish;
 end

endmodule


module park(front,back,slot,clk,start,pswd,vn);
parameter n=4;
parameter PASSWORD= 4'b1010;
parameter CLOSE=1'b0 , OPEN= 1'b1;

output reg front,back;
output reg [3:0] slot;
input start,clk;
input [n-1:0] pswd,vn;

reg [n-1:0] park[0:15];
reg [n-1:0] c_pswd;
reg f,b,state,gate;
reg k=0;

always @(posedge clk)
begin
state<=gate;
end

always@ (*)
begin
case (state)
 CLOSE: begin
	 
	 if(start)
	  begin
	   front= 1'b1;
	   c_pswd= pswd;
	   gate= OPEN;
	  end
	 else if(!start)
	  begin
	   front= 1'b0;
           back=1'b0;
	   slot=0;
	   c_pswd=0;
	   gate= CLOSE;
	  end
	end

  OPEN: begin
	 c_pswd=pswd;
	 if(c_pswd== PASSWORD)
	  begin
	    park[k]= vn;
	    slot= vn;
	    k= k+1;
	    back=1'b1;
	    gate= CLOSE;
	   end
	  else if(c_pswd!= PASSWORD)
	    begin
	    back=1'b0;
	    slot=0;
	    gate= OPEN;
	   end
	end
  default : gate= CLOSE;
 endcase

end

endmodule


 



